module client
import src.websocket as ws

fn placeholder() {}