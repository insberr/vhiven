module websocket

pub fn new_websocket() {
	println('New websocket created')
}