module hiven

pub fn hello() string {
    return 'Hello World'
}
