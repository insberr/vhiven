module rest
/*
import net.http

pub fn send(content string) {
	http.post_json('https://api.hiven.io/v1/rooms/$id/messages')
}
*/
pub fn test() {
	println('rest tested (not really)')
}