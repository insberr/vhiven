module rest

pub fn test() {
	println('rest tested (not really)')
}