module vhiven

pub fn hello() {
	println('Hello World!')
}